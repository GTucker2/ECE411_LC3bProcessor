module mux8 #(parameter width = 32)
(
	input [2:0] sel,
	input [width-1:0] a, b, c, d, e, f, g, h,
	output logic [width-1:0] i
);

always_comb
begin
	if (sel == 3'b000)
		i = a;
	else if (sel == 3'b001)
		i = b;
	else if (sel == 3'b010)
		i = c;
	else if (sel == 3'b011)
		i = d;
	else if (sel == 3'b100)
		i = e;
	else if (sel == 3'b101)
		i = f;
	else if (sel == 3'b110)
		i = g;
	else
		i = h;
end

endmodule : mux8